`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Univeristy of Washington
// Engineer: 
// 
// Create Date:    14:24:32 12/29/2013 
// Design Name: 
// Module Name:    fifos 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fifos(
	input 	rst,
	input		clk_25,
	input		clk_5,
	input		wr_en1,
	input		wr_en2,
	input		rd_en1,
	input		rd_en2,
	input		datain,
	input  [7:0] rxData,
	output problem,
	output wr_ack,
	output rd_ack,
	output [7:0] cmd,
	output [7:0] txData,
	output empty1,
	output empty2,
	output [10:0] wr_data_count // output [10 : 0] wr_data_count
    );
	 
//wire [7:0] cmd;
//wire [10:0] wr_data_count;

//generated by coregen. 8 bit to 8 bit fifo, independant read/write clocks.
cmd_fifo fifo1 (
  .rst(rst), // input rst
  .wr_clk(clk_25), // input wr_clk
  .rd_clk(clk_5), // input rd_clk
  .din(rxData), // input [7 : 0] din
  .wr_en(wr_en1), // input wr_en
  .rd_en(rd_en1), // input rd_en
  .wr_ack(wr_ack),
  .dout(cmd[7:0]), // output [7 : 0] dout
  .full(full1), // output full
  .empty(empty1), // output empty
  .wr_data_count(wr_data_count[10:0]) // output [10 : 0] wr_data_count
);

//generated by coregen. 1 bit to 8 bit fifo, independant read/write clocks.
//Possible modification in the future to 1 bit to 1 bit fifo, and then pad the
//uart tx bytes somewhere else. 
data_in_fifo fifo2 (
  .rst(rst), // input rst
  .wr_clk(clk_5), // input wr_clk
  .rd_clk(clk_25), // input rd_clk
  .din(datain), // input [0 : 0] din
  .wr_en(wr_en2), // input wr_en
  .rd_en(rd_en2), // input rd_en
  .valid(rd_ack),
  .dout(txData[7]), // output [7 : 0] dout
  .full(full2), // output full
  .empty(empty2) // output empty
);

assign txData[6] = txData[7];
assign txData[5:4] = txData[7:6];
assign txData[3:0] = txData[7:4];

assign problem = full1 || full2 || (empty1 && empty2); //simple logic to send out problem signal

endmodule
